module FOURTH_K_MAPS(
    input a,
    input b,
    input c,
    input d,
    output out  ); 
    xor(out,a,b,c,d);
endmodule

