module FIRST_K_MAPS(
    input a,
    input b,
    input c,
    output out  ); 
 assign out = a|b|c;
endmodule
